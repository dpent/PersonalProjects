library ieee;
use ieee.std_logic_1164.all;

entity and_gate2 is
	port(a, b: in std_logic;
		  c: out std_logic);
end and_gate2;


architecture behavioral of and_gate2 is
begin
	c<= a and b;
end behavioral;